library verilog;
use verilog.vl_types.all;
entity DivFrec_vlg_vec_tst is
end DivFrec_vlg_vec_tst;
