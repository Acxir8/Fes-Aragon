library verilog;
use verilog.vl_types.all;
entity Blink_vlg_vec_tst is
end Blink_vlg_vec_tst;
