library verilog;
use verilog.vl_types.all;
entity Conta_vlg_vec_tst is
end Conta_vlg_vec_tst;
