library verilog;
use verilog.vl_types.all;
entity Blink3_vlg_vec_tst is
end Blink3_vlg_vec_tst;
