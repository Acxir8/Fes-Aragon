library verilog;
use verilog.vl_types.all;
entity DIV_vlg_check_tst is
    port(
        periodo         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end DIV_vlg_check_tst;
