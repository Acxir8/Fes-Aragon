library verilog;
use verilog.vl_types.all;
entity Exceso3_vlg_vec_tst is
end Exceso3_vlg_vec_tst;
