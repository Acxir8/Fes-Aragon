library verilog;
use verilog.vl_types.all;
entity Exceso3_vlg_check_tst is
    port(
        w               : in     vl_logic;
        x               : in     vl_logic;
        y               : in     vl_logic;
        z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Exceso3_vlg_check_tst;
