library verilog;
use verilog.vl_types.all;
entity luces_vlg_vec_tst is
end luces_vlg_vec_tst;
