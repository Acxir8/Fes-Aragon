library verilog;
use verilog.vl_types.all;
entity myAND_vlg_vec_tst is
end myAND_vlg_vec_tst;
