library verilog;
use verilog.vl_types.all;
entity DIV_vlg_vec_tst is
end DIV_vlg_vec_tst;
