library verilog;
use verilog.vl_types.all;
entity semaforo_vlg_vec_tst is
end semaforo_vlg_vec_tst;
