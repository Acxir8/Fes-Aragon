module myNOT(input a, output z);
	assign z = ~a;
endmodule
