library verilog;
use verilog.vl_types.all;
entity Blink2_vlg_vec_tst is
end Blink2_vlg_vec_tst;
