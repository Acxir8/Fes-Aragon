library verilog;
use verilog.vl_types.all;
entity CarritoMueve_vlg_vec_tst is
end CarritoMueve_vlg_vec_tst;
